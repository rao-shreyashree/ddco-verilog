// This module implements a one-input NOT gate

module not_gate
(
    input a,
    output y
);

    assign y = !a;

endmodule